CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
100 150 30 150 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.499203 0.500000
344 176 1532 488
76546066 256
0
6 Title:
5 Name:
0
0
0
23
13 Logic Switch~
5 123 486 0 1 11
0 4
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 CP
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6357 0 0
2
43382.8 1
0
13 Logic Switch~
5 123 522 0 10 11
0 3 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-7 -16 7 -8
2 PL
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
319 0 0
2
43382.8 0
0
13 Logic Switch~
5 108 348 0 1 11
0 6
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 D8
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3976 0 0
2
43382.8 7
0
13 Logic Switch~
5 297 348 0 10 11
0 13 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
3 D15
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
7634 0 0
2
43382.8 6
0
13 Logic Switch~
5 270 348 0 1 11
0 12
0
0 0 21360 270
2 0V
-6 -21 8 -13
3 D14
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
523 0 0
2
43382.8 5
0
13 Logic Switch~
5 243 348 0 1 11
0 11
0
0 0 21360 270
2 0V
-6 -21 8 -13
3 D13
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6748 0 0
2
43382.8 4
0
13 Logic Switch~
5 216 348 0 1 11
0 10
0
0 0 21360 270
2 0V
-6 -21 8 -13
3 D12
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6901 0 0
2
43382.8 3
0
13 Logic Switch~
5 189 348 0 1 11
0 9
0
0 0 21360 270
2 0V
-6 -21 8 -13
3 D11
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
842 0 0
2
43382.8 2
0
13 Logic Switch~
5 162 348 0 1 11
0 8
0
0 0 21360 270
2 0V
-6 -21 8 -13
3 D10
-9 -31 12 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3277 0 0
2
43382.8 1
0
13 Logic Switch~
5 135 348 0 1 11
0 7
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 D9
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
4212 0 0
2
43382.8 0
0
13 Logic Switch~
5 135 186 0 10 11
0 17 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 D1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
4720 0 0
2
43382.8 6
0
13 Logic Switch~
5 162 186 0 10 11
0 18 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 D2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
5551 0 0
2
43382.8 5
0
13 Logic Switch~
5 189 186 0 10 11
0 19 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 D3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
6986 0 0
2
43382.8 4
0
13 Logic Switch~
5 216 186 0 10 11
0 20 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 D4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
8745 0 0
2
43382.8 3
0
13 Logic Switch~
5 243 186 0 10 11
0 21 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 D5
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
9592 0 0
2
43382.8 2
0
13 Logic Switch~
5 270 186 0 10 11
0 22 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 D6
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
8748 0 0
2
43382.8 1
0
13 Logic Switch~
5 297 186 0 10 11
0 23 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 D7
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
7168 0 0
2
43382.8 0
0
13 Logic Switch~
5 108 186 0 10 11
0 16 0 0 0 0 0 0 0 0
1
0
0 0 21360 270
2 5V
-6 -21 8 -13
2 D0
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -2 0
1 V
631 0 0
2
43382.8 0
0
14 Logic Display~
6 486 414 0 1 2
10 14
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9466 0 0
2
43382.8 0
0
7 74LS165
97 374 405 0 14 29
0 13 12 11 10 9 8 7 6 15
3 2 4 24 14
0
0 0 13040 0
7 74LS165
-24 -60 25 -52
2 U2
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 6 5 4 3 14 13 12 11 10
1 15 2 7 9 6 5 4 3 14
13 12 11 10 1 15 2 7 9 0
65 0 0 512 1 1 0 0
1 U
3266 0 0
2
43382.8 2
0
7 Ground~
168 423 414 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7693 0 0
2
43382.8 0
0
7 Ground~
168 423 252 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
3723 0 0
2
43382.8 0
0
7 74LS165
97 374 243 0 14 29
0 23 22 21 20 19 18 17 16 2
3 2 4 25 15
0
0 0 15088 0
7 74LS165
-24 -60 25 -52
2 U1
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 6 5 4 3 14 13 12 11 10
1 15 2 7 9 6 5 4 3 14
13 12 11 10 1 15 2 7 9 42
65 0 0 512 1 1 0 0
1 U
3440 0 0
2
43382.8 0
0
42
9 0 2 0 0 8192 0 23 0 0 26 3
406 207
423 207
423 225
0 1 3 0 0 8320 0 0 2 24 0 3
460 375
460 522
135 522
0 1 4 0 0 8320 0 0 1 21 0 3
441 396
441 486
135 486
0 0 5 0 0 0 0 0 0 0 0 2
288 297
288 297
8 0 6 0 0 4224 0 20 0 0 20 2
342 441
108 441
7 0 7 0 0 4224 0 20 0 0 14 2
342 432
135 432
6 0 8 0 0 4224 0 20 0 0 15 2
342 423
162 423
5 0 9 0 0 4224 0 20 0 0 13 2
342 414
189 414
4 0 10 0 0 4224 0 20 0 0 16 2
342 405
216 405
3 0 11 0 0 4224 0 20 0 0 17 2
342 396
243 396
2 0 12 0 0 4096 0 20 0 0 18 2
342 387
270 387
1 0 13 0 0 4096 0 20 0 0 19 2
342 378
297 378
1 0 9 0 0 0 0 8 0 0 0 2
189 360
189 448
1 0 7 0 0 0 0 10 0 0 0 2
135 360
135 451
1 0 8 0 0 0 0 9 0 0 0 2
162 360
162 450
1 0 10 0 0 0 0 7 0 0 0 2
216 360
216 453
1 0 11 0 0 0 0 6 0 0 0 2
243 360
243 453
1 0 12 0 0 4224 0 5 0 0 0 2
270 360
270 456
1 0 13 0 0 4224 0 4 0 0 0 2
297 360
297 455
1 0 6 0 0 0 0 3 0 0 0 2
108 360
108 453
12 12 4 0 0 0 0 23 20 0 0 4
406 234
441 234
441 396
406 396
1 14 14 0 0 8320 0 19 20 0 0 3
486 432
486 441
406 441
14 9 15 0 0 8320 0 23 20 0 0 4
406 279
414 279
414 369
406 369
10 10 3 0 0 0 0 23 20 0 0 4
412 216
460 216
460 378
412 378
1 11 2 0 0 4224 0 21 20 0 0 3
423 408
423 387
412 387
1 11 2 0 0 0 0 22 23 0 0 3
423 246
423 225
412 225
8 0 16 0 0 4224 0 23 0 0 42 2
342 279
108 279
7 0 17 0 0 4224 0 23 0 0 36 2
342 270
135 270
6 0 18 0 0 4224 0 23 0 0 37 2
342 261
162 261
5 0 19 0 0 4224 0 23 0 0 35 2
342 252
189 252
4 0 20 0 0 4224 0 23 0 0 38 2
342 243
216 243
3 0 21 0 0 4224 0 23 0 0 39 2
342 234
243 234
2 0 22 0 0 4096 0 23 0 0 40 2
342 225
270 225
1 0 23 0 0 4096 0 23 0 0 41 2
342 216
297 216
1 0 19 0 0 0 0 13 0 0 0 2
189 198
189 286
1 0 17 0 0 0 0 11 0 0 0 2
135 198
135 289
1 0 18 0 0 0 0 12 0 0 0 2
162 198
162 288
1 0 20 0 0 128 0 14 0 0 0 2
216 198
216 291
1 0 21 0 0 128 0 15 0 0 0 2
243 198
243 291
1 0 22 0 0 4224 0 16 0 0 0 2
270 198
270 294
1 0 23 0 0 4224 0 17 0 0 0 2
297 198
297 293
1 0 16 0 0 0 0 18 0 0 0 2
108 198
108 291
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
